library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package BresenhamPackage is
  -- definieer hier de functie AbsVal om de absolute waarde te
  -- berekenen van een integer
end BresenhamPackage;

package body BresenhamPackage is
end BresenhamPackage;
